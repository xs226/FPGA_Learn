module seg_led (
	clk,
	rst_n,
	segment,
	segsel
);

input clk ;
input rst_n;

output[7:0] segment;
output[7:0] segsel;
reg[7:0] segment;
reg[7:0] segsel;

parameter DATA0   = 8'b00000011  ;
parameter DATA1   = 8'b11110011  ;
parameter DATA2   = 8'b00100101  ;
parameter DATA3   = 8'b00001101  ;
parameter DATA4   = 8'b10011001  ;
parameter DATA5   = 8'b01001001  ;
parameter DATA6   = 8'b01000001  ;
parameter DATA7   = 8'b00011111  ;
parameter DATA8   = 8'b00000001  ;
parameter DATA9   = 8'b00001001  ;

parameter TIME_1s = 50_000_000 ;
reg[23:0] cnt_1s;

always @(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        cnt_1s <= 0;
    end
    else begin
        if(cnt_1s==TIME_1s-1) cnt_1s <= 0;
        else cnt_1s <= cnt_1s + 1;
    end
end

always@(posedge clk or negedge rst_n)begin
    if(rst_n==1'b0)begin
        dis_value<=0;
    end
    else if(count_20us==cnt_thd-1 && cnt_1s==TIME_1s-1 ) begin
		if(dis_value==7) dis_value<=0;
		else dis_value<=dis_value+1;
    end
end


reg[3:0] shi_s,shi_g,fen_s,fen_g,miao_s,miao_g;

always@(posedge clk or negedge rst_n)begin
    if(rst_n==1'b0)begin
        miao_g<=0;
    end
    else if(cnt_1s==TIME_1s-1) begin
        if( miao_g==9 ) miao_g<=0;
		else miao_g<=miao_g+1；
end
always@(posedge clk or negedge rst_n)begin
    if(rst_n==1'b0)begin
        miao_s<=0;
    end
    else if( miao_g==9 && cnt_1s==TIME_1s-1) begin
        if( miao_s==5 ) miao_s<=0;
		else miao_s<=miao_s+1；
end


always@(posedge clk or negedge rst_n)begin
    if(rst_n==1'b0)begin
        fen_g<=0;
    end
    else if(miao_s==5 && miao_g==9 && cnt_1s==TIME_1s-1) begin
        if( fen_g==9 ) fen_g<=0;
		else fen_g<=fen_g+1；
end
always@(posedge clk or negedge rst_n)begin
    if(rst_n==1'b0)begin
        fen_s<=0;
    end
    else if( fen_g==9 && miao_s==5 && miao_g==9 && cnt_1s==TIME_1s-1) begin
        if( fen_s==5 ) fen_s<=0;
		else fen_s<=fen_s+1；
end

always@(posedge clk or negedge rst_n)begin
    if(rst_n==1'b0)begin
        shi_g<=0;
    end
    else if(miao_s==5 && miao_g==9 && cnt_1s==TIME_1s-1) begin
		if( (shi_s<2 && shi_g==9)||(shi_s==2 && shi_g==3) shi_g<=0;
		else shi_g<=shi_g+1；
end
always@(posedge clk or negedge rst_n)begin
    if(rst_n==1'b0)begin
        shi_s<=0;
    end
    else if(shi_s<2 &&fen_g==9 && miao_s==5 && miao_g==9 && cnt_1s==TIME_1s-1)
	
	begin
        if( shi_s==2 ) fen_s<=0;
		else shi_s<=shi_s+1；
end



parameter TIME_20us = 1000 ;
reg[9:0] cnt_20us;
reg[5:0] dis_value;

always @(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        cnt_20us <= 0;
    end
    else begin
        if(cnt_20us==TIME_20us-1) cnt_20us <= 0;
        else cnt_20us <= cnt_20us + 1;
    end
end

always@(posedge clk or negedge rst_n)begin
    if(rst_n==1'b0)begin
        segsel<=8'hfe;
    end
    else if(cnt_20us==TIME_20us-1) begin
		segsel<={segsel[6:0],segsel[7]};		
    end
end

always@(*)begin
	case( dis_value )
        0:  segment <= DATA0      ;
        1:  segment <= DATA1      ;
        2:  segment <= DATA2      ;
        3:  segment <= DATA3      ;
        4:  segment <= DATA4      ;
        5:  segment <= DATA5      ;
        6:  segment <= DATA6      ;
        7:  segment <= DATA7      ;
        8:  segment <= DATA8      ;
        9:  segment <= DATA9      ;
        default:segment <= 8'hff  ;
    endcase
end


endmodule





















